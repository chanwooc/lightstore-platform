// needed by ControllerTypes.bsv
